library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity choose32 is
port(
	
	input	: in std_logic_vector(8 downto 0);
	outputA, outputB : out std_logic_vector(4 downto 0));
	
end choose32;

architecture behavioral of choose32 is
begin

	process(input)
	begin
		
		case input is
		
			-- 0,1 -> 0,31
			when "000000000" =>
				outputA <= "00000";
				outputB <= "00001";
			when "000000001" =>
				outputA <= "00000";
				outputB <= "00010";
			when "000000010" =>
				outputA <= "00000";
				outputB <= "00011";
			when "000000011" =>
				outputA <= "00000";
				outputB <= "00100";
			when "000000100" =>
				outputA <= "00000";
				outputB <= "00101";
			when "000000101" =>
				outputA <= "00000";
				outputB <= "00110";
			when "000000110" =>
				outputA <= "00000";
				outputB <= "00111";
			when "000000111" =>
				outputA <= "00000";
				outputB <= "01000";
			when "000001000" =>
				outputA <= "00000";
				outputB <= "01001";
			when "000001001" =>
				outputA <= "00000";
				outputB <= "01010";
			when "000001010" =>
				outputA <= "00000";
				outputB <= "01011";
			when "000001011" =>
				outputA <= "00000";
				outputB <= "01100";
			when "000001100" =>
				outputA <= "00000";
				outputB <= "01101";
			when "000001101" =>
				outputA <= "00000";
				outputB <= "01110";
			when "000001110" =>
				outputA <= "00000";
				outputB <= "01111";
			when "000001111" =>
				outputA <= "00000";
				outputB <= "10000";
			when "000010000" =>
				outputA <= "00000";
				outputB <= "10001";
			when "000010001" =>
				outputA <= "00000";
				outputB <= "10010";
			when "000010010" =>
				outputA <= "00000";
				outputB <= "10011";
			when "000010011" =>
				outputA <= "00000";
				outputB <= "10100";
			when "000010100" =>
				outputA <= "00000";
				outputB <= "10101";
			when "000010101" =>
				outputA <= "00000";
				outputB <= "10110";
			when "000010110" =>
				outputA <= "00000";
				outputB <= "10111";
			when "000010111" =>
				outputA <= "00000";
				outputB <= "11000";
			when "000011000" =>
				outputA <= "00000";
				outputB <= "11001";
			when "000011001" =>
				outputA <= "00000";
				outputB <= "11010";
			when "000011010" =>
				outputA <= "00000";
				outputB <= "11011";
			when "000011011" =>
				outputA <= "00000";
				outputB <= "11100";
			when "000011100" =>
				outputA <= "00000";
				outputB <= "11101";
			when "000011101" =>
				outputA <= "00000";
				outputB <= "11110";
			when "000011110" =>
				outputA <= "00000";
				outputB <= "11111";
				
			--1,2 -> 1,31
			when "000011111" =>
				outputA <= "00001";
				outputB <= "00010";
			when "000100000" =>
				outputA <= "00001";
				outputB <= "00011";
			when "000100001" =>
				outputA <= "00001";
				outputB <= "00100";
			when "000100010" =>
				outputA <= "00001";
				outputB <= "00101";
			when "000100011" =>
				outputA <= "00001";
				outputB <= "00110";
			when "000100100" =>
				outputA <= "00001";
				outputB <= "00111";
			when "000100101" =>
				outputA <= "00001";
				outputB <= "01000";
			when "000100110" =>
				outputA <= "00001";
				outputB <= "01001";
			when "000100111" =>
				outputA <= "00001";
				outputB <= "01010";
			when "000101000" =>
				outputA <= "00001";
				outputB <= "01011";
			when "000101001" =>
				outputA <= "00001";
				outputB <= "01100";
			when "000101010" =>
				outputA <= "00001";
				outputB <= "01101";
			when "000101011" =>
				outputA <= "00001";
				outputB <= "01110";
			when "000101100" =>
				outputA <= "00001";
				outputB <= "01111";
			when "000101101" =>
				outputA <= "00001";
				outputB <= "10000";
			when "000101110" =>
				outputA <= "00001";
				outputB <= "10001";
			when "000101111" =>
				outputA <= "00001";
				outputB <= "10010";
			when "000110000" =>
				outputA <= "00001";
				outputB <= "10011";
			when "000110001" =>
				outputA <= "00001";
				outputB <= "10100";
			when "000110010" =>
				outputA <= "00001";
				outputB <= "10101";
			when "000110011" =>
				outputA <= "00001";
				outputB <= "10110";
			when "000110100" =>
				outputA <= "00001";
				outputB <= "10111";
			when "000110101" =>
				outputA <= "00001";
				outputB <= "11000";
			when "000110110" =>
				outputA <= "00001";
				outputB <= "11001";
			when "000110111" =>
				outputA <= "00001";
				outputB <= "11010";
			when "000111000" =>
				outputA <= "00001";
				outputB <= "11011";
			when "000111001" =>
				outputA <= "00001";
				outputB <= "11100";
			when "000111010" =>
				outputA <= "00001";
				outputB <= "11101";
			when "000111011" =>
				outputA <= "00001";
				outputB <= "11110";
			when "000111100" =>
				outputA <= "00001";
				outputB <= "11111";
				
			-- 2,3 -> 2,31	
			when "000111101" =>
				outputA <= "00010";
				outputB <= "00011";
			when "000111110" =>
				outputA <= "00010";
				outputB <= "00100";
			when "000111111" =>	
				outputA <= "00010";
				outputB <= "00101";					
			when "001000000" =>
				outputA <= "00010";
				outputB <= "00110";
			when "001000001" =>
				outputA <= "00010";
				outputB <= "00111";
			when "001000010" =>
				outputA <= "00010";
				outputB <= "01000";
			when "001000011" =>
				outputA <= "00010";
				outputB <= "01001";
			when "001000100" =>
				outputA <= "00010";
				outputB <= "01010";
			when "001000101" =>
				outputA <= "00010";
				outputB <= "01011";
			when "001000110" =>
				outputA <= "00010";
				outputB <= "01100";
			when "001000111" =>
				outputA <= "00010";
				outputB <= "01101";
			when "001001000" =>
				outputA <= "00010";
				outputB <= "01110";
			when "001001001" =>
				outputA <= "00010";
				outputB <= "01111";
			when "001001010" =>
				outputA <= "00010";
				outputB <= "10000";
			when "001001011" =>
				outputA <= "00010";
				outputB <= "10001";
			when "001001100" =>
				outputA <= "00010";
				outputB <= "10010";
			when "001001101" =>
				outputA <= "00010";
				outputB <= "10011";
			when "001001110" =>
				outputA <= "00010";
				outputB <= "10100";
			when "001001111" =>
				outputA <= "00010";
				outputB <= "10101";
			when "001010000" =>
				outputA <= "00010";
				outputB <= "10110";
			when "001010001" =>
				outputA <= "00010";
				outputB <= "10111";
			when "001010010" =>
				outputA <= "00010";
				outputB <= "11000";
			when "001010011" =>
				outputA <= "00010";
				outputB <= "11001";
			when "001010100" =>
				outputA <= "00010";
				outputB <= "11010";
			when "001010101" =>
				outputA <= "00010";
				outputB <= "11011";
			when "001010110" =>
				outputA <= "00010";
				outputB <= "11100";
			when "001010111" =>
				outputA <= "00010";
				outputB <= "11101";
			when "001011000" =>
				outputA <= "00010";
				outputB <= "11110";
			when "001011001" =>
				outputA <= "00010";
				outputB <= "11111";
				
			-- 3,4 -> 3,31
			when "001011010" =>
				outputA <= "00011";
				outputB <= "00100";
			when "001011011" =>
				outputA <= "00011";
				outputB <= "00101";
			when "001011100" =>
				outputA <= "00011";
				outputB <= "00110";
			when "001011101" =>
				outputA <= "00011";
				outputB <= "00111";
			when "001011110" =>
				outputA <= "00011";
				outputB <= "01000";
			when "001011111" =>
				outputA <= "00011";
				outputB <= "01001";
			when "001100000" =>
				outputA <= "00011";
				outputB <= "01010";
			when "001100001" =>
				outputA <= "00011";
				outputB <= "01011";
			when "001100010" =>
				outputA <= "00011";
				outputB <= "01100";
			when "001100011" =>
				outputA <= "00011";
				outputB <= "01101";
			when "001100100" =>
				outputA <= "00011";
				outputB <= "01110";
			when "001100101" =>
				outputA <= "00011";
				outputB <= "01111";
			when "001100110" =>
				outputA <= "00011";
				outputB <= "10000";
			when "001100111" =>
				outputA <= "00011";
				outputB <= "10001";
			when "001101000" =>
				outputA <= "00011";
				outputB <= "10010";
			when "001101001" =>
				outputA <= "00011";
				outputB <= "10011";
			when "001101010" =>
				outputA <= "00011";
				outputB <= "10100";
			when "001101011" =>
				outputA <= "00011";
				outputB <= "10101";
			when "001101100" =>
				outputA <= "00011";
				outputB <= "10110";
			when "001101101" =>
				outputA <= "00011";
				outputB <= "10111";
			when "001101110" =>
				outputA <= "00011";
				outputB <= "11000";
			when "001101111" =>
				outputA <= "00011";
				outputB <= "11001";
			when "001110000" =>
				outputA <= "00011";
				outputB <= "11010";
			when "001110001" =>
				outputA <= "00011";
				outputB <= "11011";
			when "001110010" =>
				outputA <= "00011";
				outputB <= "11100";
			when "001110011" =>
				outputA <= "00011";
				outputB <= "11101";
			when "001110100" =>
				outputA <= "00011";
				outputB <= "11110";
			when "001110101" =>
				outputA <= "00011";
				outputB <= "11111";
	
			--4,5 -> 4, 31
			when "001110110" =>
				outputA <= "00100";
				outputB <= "00101";
			when "001110111" =>
				outputA <= "00100";
				outputB <= "00110";
			when "001111000" =>
				outputA <= "00100";
				outputB <= "00111";
			when "001111001" =>
				outputA <= "00100";
				outputB <= "01000";
			when "001111010" =>
				outputA <= "00100";
				outputB <= "01001";
			when "001111011" =>
				outputA <= "00100";
				outputB <= "01010";
			when "001111100" =>
				outputA <= "00100";
				outputB <= "01011";
			when "001111101" =>
				outputA <= "00100";
				outputB <= "01100";
			when "001111110" =>
				outputA <= "00100";
				outputB <= "01101";
			when "001111111" =>	
				outputA <= "00100";
				outputB <= "01110";		
			when "010000000" =>
				outputA <= "00100";
				outputB <= "01111";
			when "010000001" =>
				outputA <= "00100";
				outputB <= "10000";
			when "010000010" =>
				outputA <= "00100";
				outputB <= "10001";
			when "010000011" =>
				outputA <= "00100";
				outputB <= "10010";
			when "010000100" =>
				outputA <= "00100";
				outputB <= "10011";
			when "010000101" =>
				outputA <= "00100";
				outputB <= "10100";
			when "010000110" =>
				outputA <= "00100";
				outputB <= "10101";
			when "010000111" =>
				outputA <= "00100";
				outputB <= "10110";
			when "010001000" =>
				outputA <= "00100";
				outputB <= "10111";
			when "010001001" =>
				outputA <= "00100";
				outputB <= "11000";
			when "010001010" =>
				outputA <= "00100";
				outputB <= "11001";
			when "010001011" =>
				outputA <= "00100";
				outputB <= "11010";
			when "010001100" =>
				outputA <= "00100";
				outputB <= "11011";
			when "010001101" =>
				outputA <= "00100";
				outputB <= "11100";
			when "010001110" =>
				outputA <= "00100";
				outputB <= "11101";
			when "010001111" =>
				outputA <= "00100";
				outputB <= "11110";
			when "010010000" =>
				outputA <= "00100";
				outputB <= "11111";
				
			--5,6 -> 5,31	
			when "010010001" =>
				outputA <= "00101";
				outputB <= "00110";
			when "010010010" =>
				outputA <= "00101";
				outputB <= "00111";
			when "010010011" =>
				outputA <= "00101";
				outputB <= "01000";
			when "010010100" =>
				outputA <= "00101";
				outputB <= "01001";
			when "010010101" =>
				outputA <= "00101";
				outputB <= "01010";
			when "010010110" =>
				outputA <= "00101";
				outputB <= "01011";
			when "010010111" =>
				outputA <= "00101";
				outputB <= "01100";
			when "010011000" =>
				outputA <= "00101";
				outputB <= "01101";
			when "010011001" =>
				outputA <= "00101";
				outputB <= "01110";
			when "010011010" =>
				outputA <= "00101";
				outputB <= "01111";
			when "010011011" =>
				outputA <= "00101";
				outputB <= "10000";
			when "010011100" =>
				outputA <= "00101";
				outputB <= "10001";
			when "010011101" =>
				outputA <= "00101";
				outputB <= "10010";
			when "010011110" =>
				outputA <= "00101";
				outputB <= "10011";
			when "010011111" =>
				outputA <= "00101";
				outputB <= "10100";
			when "010100000" =>
				outputA <= "00101";
				outputB <= "10101";
			when "010100001" =>
				outputA <= "00101";
				outputB <= "10110";
			when "010100010" =>
				outputA <= "00101";
				outputB <= "10111";
			when "010100011" =>
				outputA <= "00101";
				outputB <= "11000";
			when "010100100" =>
				outputA <= "00101";
				outputB <= "11001";
			when "010100101" =>
				outputA <= "00101";
				outputB <= "11010";
			when "010100110" =>
				outputA <= "00101";
				outputB <= "11011";
			when "010100111" =>
				outputA <= "00101";
				outputB <= "11100";
			when "010101000" =>
				outputA <= "00101";
				outputB <= "11101";
			when "010101001" =>
				outputA <= "00101";
				outputB <= "11110";
			when "010101010" =>
				outputA <= "00101";
				outputB <= "11111";
				
			-- 6,7 -> 6,31	
			when "010101011" =>
				outputA <= "00110";
				outputB <= "00111";
			when "010101100" =>
				outputA <= "00110";
				outputB <= "01000";
			when "010101101" =>
				outputA <= "00110";
				outputB <= "01001";
			when "010101110" =>
				outputA <= "00110";
				outputB <= "01010";
			when "010101111" =>
				outputA <= "00110";
				outputB <= "01011";
			when "010110000" =>
				outputA <= "00110";
				outputB <= "01100";
			when "010110001" =>
				outputA <= "00110";
				outputB <= "01101";
			when "010110010" =>
				outputA <= "00110";
				outputB <= "01110";
			when "010110011" =>
				outputA <= "00110";
				outputB <= "01111";
			when "010110100" =>
				outputA <= "00110";
				outputB <= "10000";
			when "010110101" =>
				outputA <= "00110";
				outputB <= "10001";
			when "010110110" =>
				outputA <= "00110";
				outputB <= "10010";
			when "010110111" =>
				outputA <= "00110";
				outputB <= "10011";
			when "010111000" =>
				outputA <= "00110";
				outputB <= "10100";
			when "010111001" =>
				outputA <= "00110";
				outputB <= "10101";
			when "010111010" =>
				outputA <= "00110";
				outputB <= "10110";
			when "010111011" =>
				outputA <= "00110";
				outputB <= "10111";
			when "010111100" =>
				outputA <= "00110";
				outputB <= "11000";
			when "010111101" =>
				outputA <= "00110";
				outputB <= "11001";
			when "010111110" =>
				outputA <= "00110";
				outputB <= "11010";
			when "010111111" =>	
				outputA <= "00110";
				outputB <= "11011";					
			when "011000000" =>
				outputA <= "00110";
				outputB <= "11100";
			when "011000001" =>
				outputA <= "00110";
				outputB <= "11101";
			when "011000010" =>
				outputA <= "00110";
				outputB <= "11110";
			when "011000011" =>
				outputA <= "00110";
				outputB <= "11111";
				
			--7,8 -> 7,31	
			when "011000100" =>
				outputA <= "00111";
				outputB <= "01000";
			when "011000101" =>
				outputA <= "00111";
				outputB <= "01001";
			when "011000110" =>
				outputA <= "00111";
				outputB <= "01010";
			when "011000111" =>
				outputA <= "00111";
				outputB <= "01011";
			when "011001000" =>
				outputA <= "00111";
				outputB <= "01100";
			when "011001001" =>
				outputA <= "00111";
				outputB <= "01101";
			when "011001010" =>
				outputA <= "00111";
				outputB <= "01110";
			when "011001011" =>
				outputA <= "00111";
				outputB <= "01111";
			when "011001100" =>
				outputA <= "00111";
				outputB <= "10000";
			when "011001101" =>
				outputA <= "00111";
				outputB <= "10001";
			when "011001110" =>
				outputA <= "00111";
				outputB <= "10010";
			when "011001111" =>
				outputA <= "00111";
				outputB <= "10011";
			when "011010000" =>
				outputA <= "00111";
				outputB <= "10100";
			when "011010001" =>
				outputA <= "00111";
				outputB <= "10101";
			when "011010010" =>
				outputA <= "00111";
				outputB <= "10110";
			when "011010011" =>
				outputA <= "00111";
				outputB <= "10111";
			when "011010100" =>
				outputA <= "00111";
				outputB <= "11000";
			when "011010101" =>
				outputA <= "00111";
				outputB <= "11001";
			when "011010110" =>
				outputA <= "00111";
				outputB <= "11010";
			when "011010111" =>
				outputA <= "00111";
				outputB <= "11011";
			when "011011000" =>
				outputA <= "00111";
				outputB <= "11100";
			when "011011001" =>
				outputA <= "00111";
				outputB <= "11101";
			when "011011010" =>
				outputA <= "00111";
				outputB <= "11110";
			when "011011011" =>
				outputA <= "00111";
				outputB <= "11111";
				
			--8,9 -> 8,31	
			when "011011100" =>
				outputA <= "01000";
				outputB <= "01001";
			when "011011101" =>
				outputA <= "01000";
				outputB <= "01010";
			when "011011110" =>
				outputA <= "01000";
				outputB <= "01011";
			when "011011111" =>
				outputA <= "01000";
				outputB <= "01100";
			when "011100000" =>
				outputA <= "01000";
				outputB <= "01101";
			when "011100001" =>
				outputA <= "01000";
				outputB <= "01110";
			when "011100010" =>
				outputA <= "01000";
				outputB <= "01111";
			when "011100011" =>
				outputA <= "01000";
				outputB <= "10000";
			when "011100100" =>
				outputA <= "01000";
				outputB <= "10001";
			when "011100101" =>
				outputA <= "01000";
				outputB <= "10010";
			when "011100110" =>
				outputA <= "01000";
				outputB <= "10011";
			when "011100111" =>
				outputA <= "01000";
				outputB <= "10100";
			when "011101000" =>
				outputA <= "01000";
				outputB <= "10101";
			when "011101001" =>
				outputA <= "01000";
				outputB <= "10110";
			when "011101010" =>
				outputA <= "01000";
				outputB <= "10111";
			when "011101011" =>
				outputA <= "01000";
				outputB <= "11000";
			when "011101100" =>
				outputA <= "01000";
				outputB <= "11001";
			when "011101101" =>
				outputA <= "01000";
				outputB <= "11010";
			when "011101110" =>
				outputA <= "01000";
				outputB <= "11011";
			when "011101111" =>
				outputA <= "01000";
				outputB <= "11100";
			when "011110000" =>
				outputA <= "01000";
				outputB <= "11101";
			when "011110001" =>
				outputA <= "01000";
				outputB <= "11110";
			when "011110010" =>
				outputA <= "01000";
				outputB <= "11111";
				
			--9,10 -> 9,31	
			when "011110011" =>
				outputA <= "01001";
				outputB <= "01010";
			when "011110100" =>
				outputA <= "01001";
				outputB <= "01011";
			when "011110101" =>
				outputA <= "01001";
				outputB <= "01100";
			when "011110110" =>
				outputA <= "01001";
				outputB <= "01101";
			when "011110111" =>
				outputA <= "01001";
				outputB <= "01110";
			when "011111000" =>
				outputA <= "01001";
				outputB <= "01111";
			when "011111001" =>
				outputA <= "01001";
				outputB <= "10000";
			when "011111010" =>
				outputA <= "01001";
				outputB <= "10001";
			when "011111011" =>
				outputA <= "01001";
				outputB <= "10010";
			when "011111100" =>
				outputA <= "01001";
				outputB <= "10011";
			when "011111101" =>
				outputA <= "01001";
				outputB <= "10100";
			when "011111110" =>
				outputA <= "01001";
				outputB <= "10101";
			when "011111111" =>
				outputA <= "01001";
				outputB <= "10110";
			when "100000000" =>
				outputA <= "01001";
				outputB <= "10111";
			when "100000001" =>
				outputA <= "01001";
				outputB <= "11000";
			when "100000010" =>
				outputA <= "01001";
				outputB <= "11001";
			when "100000011" =>
				outputA <= "01001";
				outputB <= "11010";
			when "100000100" =>
				outputA <= "01001";
				outputB <= "11011";
			when "100000101" =>
				outputA <= "01001";
				outputB <= "11100";
			when "100000110" =>
				outputA <= "01001";
				outputB <= "11101";
			when "100000111" =>
				outputA <= "01001";
				outputB <= "11110";
			when "100001000" =>
				outputA <= "01001";
				outputB <= "11111";
				
			--10,11 -> 10,31	
			when "100001001" =>
				outputA <= "01010";
				outputB <= "01011";
			when "100001010" =>
				outputA <= "01010";
				outputB <= "01100";
			when "100001011" =>
				outputA <= "01010";
				outputB <= "01101";
			when "100001100" =>
				outputA <= "01010";
				outputB <= "01110";
			when "100001101" =>
				outputA <= "01010";
				outputB <= "01111";
			when "100001110" =>
				outputA <= "01010";
				outputB <= "10000";
			when "100001111" =>
				outputA <= "01010";
				outputB <= "10001";
			when "100010000" =>
				outputA <= "01010";
				outputB <= "10010";
			when "100010001" =>
				outputA <= "01010";
				outputB <= "10011";
			when "100010010" =>
				outputA <= "01010";
				outputB <= "10100";
			when "100010011" =>
				outputA <= "01010";
				outputB <= "10101";
			when "100010100" =>
				outputA <= "01010";
				outputB <= "10110";
			when "100010101" =>
				outputA <= "01010";
				outputB <= "10111";
			when "100010110" =>
				outputA <= "01010";
				outputB <= "11000";
			when "100010111" =>
				outputA <= "01010";
				outputB <= "11001";
			when "100011000" =>
				outputA <= "01010";
				outputB <= "11010";
			when "100011001" =>
				outputA <= "01010";
				outputB <= "11011";
			when "100011010" =>
				outputA <= "01010";
				outputB <= "11100";
			when "100011011" =>
				outputA <= "01010";
				outputB <= "11101";
			when "100011100" =>
				outputA <= "01010";
				outputB <= "11110";
			when "100011101" =>
				outputA <= "01010";
				outputB <= "11111";
				
			--11,12 -> 11,31
			when "100011110" =>
				outputA <= "01011";
				outputB <= "01100";
			when "100011111" =>
				outputA <= "01011";
				outputB <= "01101";
			when "100100000" =>
				outputA <= "01011";
				outputB <= "01110";
			when "100100001" =>
				outputA <= "01011";
				outputB <= "01111";
			when "100100010" =>
				outputA <= "01011";
				outputB <= "10000";
			when "100100011" =>
				outputA <= "01011";
				outputB <= "10001";
			when "100100100" =>
				outputA <= "01011";
				outputB <= "10010";
			when "100100101" =>
				outputA <= "01011";
				outputB <= "10011";
			when "100100110" =>
				outputA <= "01011";
				outputB <= "10100";
			when "100100111" =>
				outputA <= "01011";
				outputB <= "10101";
			when "100101000" =>
				outputA <= "01011";
				outputB <= "10110";
			when "100101001" =>
				outputA <= "01011";
				outputB <= "10111";
			when "100101010" =>
				outputA <= "01011";
				outputB <= "11000";
			when "100101011" =>
				outputA <= "01011";
				outputB <= "11001";
			when "100101100" =>
				outputA <= "01011";
				outputB <= "11010";
			when "100101101" =>
				outputA <= "01011";
				outputB <= "11011";
			when "100101110" =>
				outputA <= "01011";
				outputB <= "11100";
			when "100101111" =>
				outputA <= "01011";
				outputB <= "11101";
			when "100110000" =>
				outputA <= "01011";
				outputB <= "11110";
			when "100110001" =>
				outputA <= "01011";
				outputB <= "11111";
				
			--12,13 -> 12,31	
			when "100110010" =>
				outputA <= "01100";
				outputB <= "01101";
			when "100110011" =>
				outputA <= "01100";
				outputB <= "01110";
			when "100110100" =>
				outputA <= "01100";
				outputB <= "01111";
			when "100110101" =>
				outputA <= "01100";
				outputB <= "10000";
			when "100110110" =>
				outputA <= "01100";
				outputB <= "10001";
			when "100110111" =>
				outputA <= "01100";
				outputB <= "10010";
			when "100111000" =>
				outputA <= "01100";
				outputB <= "10011";
			when "100111001" =>
				outputA <= "01100";
				outputB <= "10100";
			when "100111010" =>
				outputA <= "01100";
				outputB <= "10101";
			when "100111011" =>
				outputA <= "01100";
				outputB <= "10110";
			when "100111100" =>
				outputA <= "01100";
				outputB <= "10111";
			when "100111101" =>
				outputA <= "01100";
				outputB <= "11000";
			when "100111110" =>
				outputA <= "01100";
				outputB <= "11001";
			when "100111111" =>	
				outputA <= "01100";
				outputB <= "11010";					
			when "101000000" =>
				outputA <= "01100";
				outputB <= "11011";
			when "101000001" =>
				outputA <= "01100";
				outputB <= "11100";
			when "101000010" =>
				outputA <= "01100";
				outputB <= "11101";
			when "101000011" =>
				outputA <= "01100";
				outputB <= "11110";
			when "101000100" =>
				outputA <= "01100";
				outputB <= "11111";
				
			--13,14 -> 13,31
			when "101000101" =>
				outputA <= "01101";
				outputB <= "01110";
			when "101000110" =>
				outputA <= "01101";
				outputB <= "01111";
			when "101000111" =>
				outputA <= "01101";
				outputB <= "10000";
			when "101001000" =>
				outputA <= "01101";
				outputB <= "10001";
			when "101001001" =>
				outputA <= "01101";
				outputB <= "10010";
			when "101001010" =>
				outputA <= "01101";
				outputB <= "10011";
			when "101001011" =>
				outputA <= "01101";
				outputB <= "10100";
			when "101001100" =>
				outputA <= "01101";
				outputB <= "10101";
			when "101001101" =>
				outputA <= "01101";
				outputB <= "10110";
			when "101001110" =>
				outputA <= "01101";
				outputB <= "10111";
			when "101001111" =>
				outputA <= "01101";
				outputB <= "11000";
			when "101010000" =>
				outputA <= "01101";
				outputB <= "11001";
			when "101010001" =>
				outputA <= "01101";
				outputB <= "11010";
			when "101010010" =>
				outputA <= "01101";
				outputB <= "11011";
			when "101010011" =>
				outputA <= "01101";
				outputB <= "11100";
			when "101010100" =>
				outputA <= "01101";
				outputB <= "11101";
			when "101010101" =>
				outputA <= "01101";
				outputB <= "11110";
			when "101010110" =>
				outputA <= "01101";
				outputB <= "11111";
				
			--14,15 -> 14,31
			when "101010111" =>
				outputA <= "01110";
				outputB <= "01111";
			when "101011000" =>
				outputA <= "01110";
				outputB <= "10000";
			when "101011001" =>
				outputA <= "01110";
				outputB <= "10001";
			when "101011010" =>
				outputA <= "01110";
				outputB <= "10010";
			when "101011011" =>
				outputA <= "01110";
				outputB <= "10011";
			when "101011100" =>
				outputA <= "01110";
				outputB <= "10100";
			when "101011101" =>
				outputA <= "01110";
				outputB <= "10101";
			when "101011110" =>
				outputA <= "01110";
				outputB <= "10110";
			when "101011111" =>
				outputA <= "01110";
				outputB <= "10111";
			when "101100000" =>
				outputA <= "01110";
				outputB <= "11000";
			when "101100001" =>
				outputA <= "01110";
				outputB <= "11001";
			when "101100010" =>
				outputA <= "01110";
				outputB <= "11010";
			when "101100011" =>
				outputA <= "01110";
				outputB <= "11011";
			when "101100100" =>
				outputA <= "01110";
				outputB <= "11100";
			when "101100101" =>
				outputA <= "01110";
				outputB <= "11101";
			when "101100110" =>
				outputA <= "01110";
				outputB <= "11110";
			when "101100111" =>
				outputA <= "01110";
				outputB <= "11111";
			
			--15,16 -> 15,31
			when "101101000" =>
				outputA <= "01111";
				outputB <= "10000";
			when "101101001" =>
				outputA <= "01111";
				outputB <= "10001";
			when "101101010" =>
				outputA <= "01111";
				outputB <= "10010";
			when "101101011" =>
				outputA <= "01111";
				outputB <= "10011";
			when "101101100" =>
				outputA <= "01111";
				outputB <= "10100";
			when "101101101" =>
				outputA <= "01111";
				outputB <= "10101";
			when "101101110" =>
				outputA <= "01111";
				outputB <= "10110";
			when "101101111" =>
				outputA <= "01111";
				outputB <= "10111";
			when "101110000" =>
				outputA <= "01111";
				outputB <= "11000";
			when "101110001" =>
				outputA <= "01111";
				outputB <= "11001";
			when "101110010" =>
				outputA <= "01111";
				outputB <= "11010";
			when "101110011" =>
				outputA <= "01111";
				outputB <= "11011";
			when "101110100" =>
				outputA <= "01111";
				outputB <= "11100";
			when "101110101" =>
				outputA <= "01111";
				outputB <= "11101";
			when "101110110" =>
				outputA <= "01111";
				outputB <= "11110";
			when "101110111" =>
				outputA <= "01111";
				outputB <= "11111";
				
			--16,17 -> 16,31
			when "101111000" =>
				outputA <= "10000";
				outputB <= "10001";
			when "101111001" =>
				outputA <= "10000";
				outputB <= "10010";
			when "101111010" =>
				outputA <= "10000";
				outputB <= "10011";
			when "101111011" =>
				outputA <= "10000";
				outputB <= "10100";
			when "101111100" =>
				outputA <= "10000";
				outputB <= "10101";
			when "101111101" =>
				outputA <= "10000";
				outputB <= "10110";
			when "101111110" =>
				outputA <= "10000";
				outputB <= "10111";
			when "101111111" =>	
				outputA <= "10000";
				outputB <= "11000";		
			when "110000000" =>
				outputA <= "10000";
				outputB <= "11001";
			when "110000001" =>
				outputA <= "10000";
				outputB <= "11010";
			when "110000010" =>
				outputA <= "10000";
				outputB <= "11011";
			when "110000011" =>
				outputA <= "10000";
				outputB <= "11100";
			when "110000100" =>
				outputA <= "10000";
				outputB <= "11101";
			when "110000101" =>
				outputA <= "10000";
				outputB <= "11110";
			when "110000110" =>
				outputA <= "10000";
				outputB <= "11111";
				
			--17,18 -> 17,31
			when "110000111" =>
				outputA <= "10001";
				outputB <= "10010";
			when "110001000" =>
				outputA <= "10001";
				outputB <= "10011";
			when "110001001" =>
				outputA <= "10001";
				outputB <= "10100";
			when "110001010" =>
				outputA <= "10001";
				outputB <= "10101";
			when "110001011" =>
				outputA <= "10001";
				outputB <= "10110";
			when "110001100" =>
				outputA <= "10001";
				outputB <= "10111";
			when "110001101" =>
				outputA <= "10001";
				outputB <= "11000";
			when "110001110" =>
				outputA <= "10001";
				outputB <= "11001";
			when "110001111" =>
				outputA <= "10001";
				outputB <= "11010";
			when "110010000" =>
				outputA <= "10001";
				outputB <= "11011";
			when "110010001" =>
				outputA <= "10001";
				outputB <= "11100";
			when "110010010" =>
				outputA <= "10001";
				outputB <= "11101";
			when "110010011" =>
				outputA <= "10001";
				outputB <= "11110";
			when "110010100" =>
				outputA <= "10001";
				outputB <= "11111";
				
			--18,19 -> 18,31
			when "110010101" =>
				outputA <= "10010";
				outputB <= "10011";
			when "110010110" =>
				outputA <= "10010";
				outputB <= "10100";
			when "110010111" =>
				outputA <= "10010";
				outputB <= "10101";
			when "110011000" =>
				outputA <= "10010";
				outputB <= "10110";
			when "110011001" =>
				outputA <= "10010";
				outputB <= "10111";
			when "110011010" =>
				outputA <= "10010";
				outputB <= "11000";
			when "110011011" =>
				outputA <= "10010";
				outputB <= "11001";
			when "110011100" =>
				outputA <= "10010";
				outputB <= "11010";
			when "110011101" =>
				outputA <= "10010";
				outputB <= "11011";
			when "110011110" =>
				outputA <= "10010";
				outputB <= "11100";
			when "110011111" =>
				outputA <= "10010";
				outputB <= "11101";
			when "110100000" =>
				outputA <= "10010";
				outputB <= "11110";
			when "110100001" =>
				outputA <= "10010";
				outputB <= "11111";
				
			--19,20 -> 19,31
			when "110100010" =>
				outputA <= "10011";
				outputB <= "10100";
			when "110100011" =>
				outputA <= "10011";
				outputB <= "10101";
			when "110100100" =>
				outputA <= "10011";
				outputB <= "10110";
			when "110100101" =>
				outputA <= "10011";
				outputB <= "10111";
			when "110100110" =>
				outputA <= "10011";
				outputB <= "11000";
			when "110100111" =>
				outputA <= "10011";
				outputB <= "11001";
			when "110101000" =>
				outputA <= "10011";
				outputB <= "11010";
			when "110101001" =>
				outputA <= "10011";
				outputB <= "11011";
			when "110101010" =>
				outputA <= "10011";
				outputB <= "11100";
			when "110101011" =>
				outputA <= "10011";
				outputB <= "11101";
			when "110101100" =>
				outputA <= "10011";
				outputB <= "11110";
			when "110101101" =>
				outputA <= "10011";
				outputB <= "11111";
				
			--20,21 -> 20,31
			when "110101110" =>
				outputA <= "10100";
				outputB <= "10101";
			when "110101111" =>
				outputA <= "10100";
				outputB <= "10110";
			when "110110000" =>
				outputA <= "10100";
				outputB <= "10111";
			when "110110001" =>
				outputA <= "10100";
				outputB <= "11000";
			when "110110010" =>
				outputA <= "10100";
				outputB <= "11001";
			when "110110011" =>
				outputA <= "10100";
				outputB <= "11010";
			when "110110100" =>
				outputA <= "10100";
				outputB <= "11011";
			when "110110101" =>
				outputA <= "10100";
				outputB <= "11100";
			when "110110110" =>
				outputA <= "10100";
				outputB <= "11101";
			when "110110111" =>
				outputA <= "10100";
				outputB <= "11110";
			when "110111000" =>
				outputA <= "10100";
				outputB <= "11111";
				
			--21,22 -> 21,31
			when "110111001" =>
				outputA <= "10101";
				outputB <= "10110";
			when "110111010" =>
				outputA <= "10101";
				outputB <= "10111";
			when "110111011" =>
				outputA <= "10101";
				outputB <= "11000";
			when "110111100" =>
				outputA <= "10101";
				outputB <= "11001";
			when "110111101" =>
				outputA <= "10101";
				outputB <= "11010";
			when "110111110" =>
				outputA <= "10101";
				outputB <= "11011";
			when "110111111" =>	
				outputA <= "10101";
				outputB <= "11100";					
			when "111000000" =>
				outputA <= "10101";
				outputB <= "11101";
			when "111000001" =>
				outputA <= "10101";
				outputB <= "11110";
			when "111000010" =>
				outputA <= "10101";
				outputB <= "11111";
				
			--22,23 -> 22,31
			when "111000011" =>
				outputA <= "10110";
				outputB <= "10111";
			when "111000100" =>
				outputA <= "10110";
				outputB <= "11000";
			when "111000101" =>
				outputA <= "10110";
				outputB <= "11001";
			when "111000110" =>
				outputA <= "10110";
				outputB <= "11010";
			when "111000111" =>
				outputA <= "10110";
				outputB <= "11011";
			when "111001000" =>
				outputA <= "10110";
				outputB <= "11100";
			when "111001001" =>
				outputA <= "10110";
				outputB <= "11101";
			when "111001010" =>
				outputA <= "10110";
				outputB <= "11110";
			when "111001011" =>
				outputA <= "10110";
				outputB <= "11111";
				
			--23,24 -> 23,31
			when "111001100" =>
				outputA <= "10111";
				outputB <= "11000";
			when "111001101" =>
				outputA <= "10111";
				outputB <= "11001";
			when "111001110" =>
				outputA <= "10111";
				outputB <= "11010";
			when "111001111" =>
				outputA <= "10111";
				outputB <= "11011";
			when "111010000" =>
				outputA <= "10111";
				outputB <= "11100";
			when "111010001" =>
				outputA <= "10111";
				outputB <= "11101";
			when "111010010" =>
				outputA <= "10111";
				outputB <= "11110";
			when "111010011" =>
				outputA <= "10111";
				outputB <= "11111";
				
			--24,25 -> 24,31
			when "111010100" =>
				outputA <= "11000";
				outputB <= "11001";
			when "111010101" =>
				outputA <= "11000";
				outputB <= "11010";
			when "111010110" =>
				outputA <= "11000";
				outputB <= "11011";
			when "111010111" =>
				outputA <= "11000";
				outputB <= "11100";
			when "111011000" =>
				outputA <= "11000";
				outputB <= "11101";
			when "111011001" =>
				outputA <= "11000";
				outputB <= "11110";
			when "111011010" =>
				outputA <= "11000";
				outputB <= "11111";
				
			--25,26 -> 25,31
			when "111011011" =>
				outputA <= "11001";
				outputB <= "11010";
			when "111011100" =>
				outputA <= "11001";
				outputB <= "11011";
			when "111011101" =>
				outputA <= "11001";
				outputB <= "11100";
			when "111011110" =>
				outputA <= "11001";
				outputB <= "11101";
			when "111011111" =>
				outputA <= "11001";
				outputB <= "11110";
			when "111100000" =>
				outputA <= "11001";
				outputB <= "11111";
				
			--26,27 -> 26,31
			when "111100001" =>
				outputA <= "11010";
				outputB <= "11011";
			when "111100010" =>
				outputA <= "11010";
				outputB <= "11100";
			when "111100011" =>
				outputA <= "11010";
				outputB <= "11101";
			when "111100100" =>
				outputA <= "11010";
				outputB <= "11110";
			when "111100101" =>
				outputA <= "11010";
				outputB <= "11111";
				
			--27,28 -> 27,31
			when "111100110" =>
				outputA <= "11011";
				outputB <= "11100";
			when "111100111" =>
				outputA <= "11011";
				outputB <= "11101";
			when "111101000" =>
				outputA <= "11011";
				outputB <= "11110";
			when "111101001" =>
				outputA <= "11011";
				outputB <= "11111";

			--28,29 -> 28,31
			when "111101010" =>
				outputA <= "11100";
				outputB <= "11101";
			when "111101011" =>
				outputA <= "11100";
				outputB <= "11110";
			when "111101100" =>
				outputA <= "11100";
				outputB <= "11111";
				
			--29,30 -> 29,31
			when "111101101" =>
				outputA <= "11101";
				outputB <= "11110";
			when "111101110" =>
				outputA <= "11101";
				outputB <= "11111";
				
			--30,31
			when "111101111" =>
				outputA <= "11110";
				outputB <= "11111";
			
			when others =>
				outputA <= "UUUUU";
				outputB <= "UUUUU";
				
		end case;
	end process;
end behavioral;